`timescale 1ns / 1ps
`default_nettype none

module keyboard_ram (
  input wire clk_in,
  input wire rst_in,
  
  output logic [7:0] scancode_out,
  
);
  
endmodule