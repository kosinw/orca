`timescale 1ns / 1ps
`default_nettype none
`include "hdl/riscv_constants.svg"

module riscv_core (
    input wire clk_in,
    input wire rst_in,

);
endmodule